module half_adder
