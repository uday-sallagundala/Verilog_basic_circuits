module half_adder_tb
